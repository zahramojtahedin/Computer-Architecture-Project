module ID(input [31:0]INSTR,WR, input [4:0]RD_ADD_IN, output [4:0]RD_ADD_OUT,RS_ADD_OUT,RT_ADD_OUT, input WE,CLK, output [31:0]IMM_OFST,RS,RT, output [2:0]OP_CAT,CMD, output UNSGN,IS_IMM,WB_EN,MEM_EN,IS_LD,IS_LDI);
parameter _non=5,_st=4,_ld=3,_br2=2,_br1=1,_ar=0;
parameter _add=0,_sub=1,_and=2,_or=3,_xor=4,_nor=5,_slt=6;
wire [5:0]OP=INSTR[31:26];
wire [4:0]RS_ADD=INSTR[25:21];
wire [4:0]RT_ADD=INSTR[20:16];
wire _unsgn=(OP==6'b100001)|(OP==6'b00011)|(OP==6'b101111)|(OP[5:1]==5'b00001)|(OP==6'b001001);
wire sgn=(!_unsgn)&INSTR[15];
assign RS_ADD_OUT=RS_ADD;
assign RT_ADD_OUT=RT_ADD;
assign UNSGN=_unsgn;
assign OP_CAT=(OP==6'b111111)?_st:(OP[5:1]==5'b10111)?_ld:(OP==6'b101000)?_br1:(OP==6'b101001)?_br2:(OP<=6'b100110)?_ar:_non;
assign WB_EN=(OP_CAT==_ld)|(OP_CAT==_ar);
assign MEM_EN=(OP_CAT==_st);
assign IS_IMM=OP[5]&&(OP_CAT!=_br1)&&(OP_CAT!=_br2)|(OP_CAT==_st);
assign IS_LD=(OP_CAT==_ld)&& !OP[0];
assign IS_LDI=(OP_CAT==_ld)&& OP[0];
assign IMM_OFST=IS_LDI?{{16{1'b0}},{INSTR[15:0]}}:{{16{sgn}},INSTR[15:0]};
assign RD_ADD_OUT=IS_IMM?RT_ADD:INSTR[15:11];
assign CMD=((OP[4:1]==4'b0000)|(OP_CAT==_ld))?_add:(OP==6'b000001)?_sub:(OP[4:0]==5'b00100)?_and:(OP[4:0]==5'b00101)?_or:(OP[4:0]==5'b00110)?_xor:(OP==6'b000111)?_nor:((OP[5:1]==5'b00100)||(OP[5:1]==5'b10001))?_slt:_add;
REG _REG (.RS_ADD(RS_ADD),.RT_ADD(RT_ADD),.RD_ADD(RD_ADD_IN),.WR(WR),.WE(WE),.CLK(CLK),.RS(RS),.RT(RT));
endmodule;