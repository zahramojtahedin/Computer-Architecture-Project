module CPU(input CLK);
wire [31:0]PC_4_MEM,PC_4_IF,INSTR_IF,INSTR_ID,PC_4_ID,WB_OUT,IMM_OFST_ID,RS_ID,RT_ID,PC_4_EX,IMM_OFST_EX,RS_EX,RT_EX,ALU_OUT_EX,ALU_OUT_MEM,RT_MEM,ALU_OUT_WB,MEM_OUT_WB,PC_4_EX_OUT,MEM_OUT_MEM;
wire IS_LDI_ID,IS_LDI_EX,IS_LDI_MEM,IS_LDI_WB,IS_LD_ID,IS_LD_EX,IS_LD_MEM,IS_LD_WB,WB_EN_WB,UNSGN_ID,IS_IMM_ID,WB_EN_ID,MEM_EN_ID,UNSGN_EX,IS_IMM_EX,WB_EN_EX,MEM_EN_EX,BRANCH_EX,BRANCH_MEM,WB_EN_MEM,MEM_EN_MEM;
wire [1:0]SELS,SELT;
wire PC_SEL,PC_WE,IS_BR_EX;
wire [2:0]OP_CAT_ID,CMD_ID,OP_CAT_EX,CMD_EX;
wire [4:0]RD_ADD_OUT_ID,RD_ADD_OUT_EX,RD_ADD_OUT_MEM,RD_ADD_OUT_WB,RS_ADD_OUT_ID,RT_ADD_OUT_ID,RS_ADD_OUT_EX,RT_ADD_OUT_EX;
wire FLUSH_BR_PRED;
IF     _IF    (.PC_4_IN(PC_4_MEM),.PC_SEL(PC_SEL),.CLK(CLK),.PC_WE(PC_WE),.PC_4_OUT(PC_4_IF),.INSTR(INSTR_IF),.IS_BR_EX(IS_BR_EX),.BRANCH_EX(BRANCH_EX),.FLUSH(FLUSH_BR_PRED));
IF_ID  _IF_ID (.RST(FLUSH_BR_PRED),.IN({PC_4_IF,INSTR_IF}),.CLK(CLK),.OUT({PC_4_ID,INSTR_ID}));
ID     _ID    (.INSTR(INSTR_ID),.WR(WB_OUT),.RD_ADD_IN(RD_ADD_OUT_WB),.RD_ADD_OUT(RD_ADD_OUT_ID),.RS_ADD_OUT(RS_ADD_OUT_ID),.RT_ADD_OUT(RT_ADD_OUT_ID),.WE(WB_EN_WB),.CLK(CLK),.IMM_OFST(IMM_OFST_ID),.RS(RS_ID),.RT(RT_ID),.OP_CAT(OP_CAT_ID),.CMD(CMD_ID),.UNSGN(UNSGN_ID),.IS_IMM(IS_IMM_ID),.WB_EN(WB_EN_ID),.MEM_EN(MEM_EN_ID),.IS_LD(IS_LD_ID),.IS_LDI(IS_LDI_ID));
ID_EX  _ID_EX (.RST(FLUSH_BR_PRED),.IN({IS_LD_ID,PC_4_ID,RD_ADD_OUT_ID,IMM_OFST_ID,RS_ID,RT_ID,OP_CAT_ID,CMD_ID,UNSGN_ID,IS_IMM_ID,WB_EN_ID,MEM_EN_ID,RS_ADD_OUT_ID,RT_ADD_OUT_ID,IS_LDI_ID}),.CLK(CLK),.OUT({IS_LD_EX,PC_4_EX,RD_ADD_OUT_EX,IMM_OFST_EX,RS_EX,RT_EX,OP_CAT_EX,CMD_EX,UNSGN_EX,IS_IMM_EX,WB_EN_EX,MEM_EN_EX,RS_ADD_OUT_EX,RT_ADD_OUT_EX,IS_LDI_EX}));
EX     _EX    (.RS(RS_EX),.RT(RT_EX),.R_MEM(ALU_OUT_MEM),.R_WB(WB_OUT),.IMM_OFST(IMM_OFST_EX),.PC_4_IN(PC_4_EX),.SELS(SELS),.SELT(SELT),.UNSGN(UNSGN_EX),.OP_CAT(OP_CAT_EX),.CMD(CMD_EX),.PC_4_OUT(PC_4_EX_OUT),.ALU_OUT(ALU_OUT_EX),.BRANCH(BRANCH_EX),.IS_BR(IS_BR_EX));
EX_MEM _EX_MEM(.RST(FLUSH_BR_PRED),.IN({IS_LD_EX,PC_4_EX_OUT,RD_ADD_OUT_EX,BRANCH_EX,ALU_OUT_EX,RT_EX,WB_EN_EX,MEM_EN_EX,IS_LDI_EX}),.CLK(CLK),.OUT({IS_LD_MEM,PC_4_MEM,RD_ADD_OUT_MEM,BRANCH_MEM,ALU_OUT_MEM,RT_MEM,WB_EN_MEM,MEM_EN_MEM,IS_LDI_MEM}));
MEM    _MEM   (.ADD(ALU_OUT_MEM[15:0]),.WR(RT_MEM),.WE(MEM_EN_MEM),.CLK(CLK),.RD(MEM_OUT_MEM));
MEM_WB _MEM_WB(.IN({IS_LD_MEM,RD_ADD_OUT_MEM,MEM_OUT_MEM,ALU_OUT_MEM,WB_EN_MEM,IS_LDI_MEM}),.CLK(CLK),.OUT({IS_LD_WB,RD_ADD_OUT_WB,MEM_OUT_WB,ALU_OUT_WB,WB_EN_WB,IS_LDI_WB}));
WB     _WB    (.MEM(MEM_OUT_WB),.ALU(ALU_OUT_WB),.SEL(IS_LD_WB),.OUT(WB_OUT));
Forwarder _Forwarder(.WB_EN_MEM(WB_EN_MEM),.WB_EN_WB(WB_EN_WB),.IS_IMM(IS_IMM_EX),.IS_LDI(IS_LDI_ID),.RS(RS_ADD_OUT_EX),.RT(RT_ADD_OUT_EX),.RD_ADD_OUT_MEM(RD_ADD_OUT_MEM),.RD_ADD_OUT_WB(RD_ADD_OUT_WB),.SELS(SELS),.SELT(SELT));
Controller _Controller(.CLK(CLK),.BRANCH(BRANCH_EX),.PC_SEL(PC_SEL),.PC_WE(PC_WE));
endmodule;
